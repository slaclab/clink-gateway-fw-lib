-------------------------------------------------------------------------------
-- Company    : SLAC National Accelerator Laboratory
-------------------------------------------------------------------------------
-- Description:
-------------------------------------------------------------------------------
-- This file is part of 'Camera link gateway'.
-- It is subject to the license terms in the LICENSE.txt file found in the
-- top-level directory of this distribution and at:
--    https://confluence.slac.stanford.edu/display/ppareg/LICENSE.html.
-- No part of 'Camera link gateway', including this file,
-- may be copied, modified, propagated, or distributed except according to
-- the terms contained in the LICENSE.txt file.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;


library surf;
use surf.StdRtlPkg.all;
use surf.AxiStreamPkg.all;
use surf.AxiLitePkg.all;
use surf.SsiPkg.all;
use surf.Pgp3Pkg.all;
use surf.ClinkPkg.all;

entity CLinkWrapper is
   generic (
      TPD_G            : time                 := 1 ns;
      CHAN_COUNT_G     : integer range 1 to 2 := 1;
      AXIL_BASE_ADDR_G : slv(31 downto 0));
   port (
      -- Clink Ports
      cbl0Half0P      : inout slv(4 downto 0);  --  2,  4,  5,  6, 3
      cbl0Half0M      : inout slv(4 downto 0);  -- 15, 17, 18, 19 16
      cbl0Half1P      : inout slv(4 downto 0);  --  8, 10, 11, 12,  9
      cbl0Half1M      : inout slv(4 downto 0);  -- 21, 23, 24, 25, 22
      cbl0SerP        : out   sl;               -- 20
      cbl0SerM        : out   sl;               -- 7
      cbl1Half0P      : inout slv(4 downto 0);  --  2,  4,  5,  6, 3
      cbl1Half0M      : inout slv(4 downto 0);  -- 15, 17, 18, 19 16
      cbl1Half1P      : inout slv(4 downto 0);  --  8, 10, 11, 12,  9
      cbl1Half1M      : inout slv(4 downto 0);  -- 21, 23, 24, 25, 22
      cbl1SerP        : out   sl;               -- 20
      cbl1SerM        : out   sl;               -- 7
      -- LEDs
      ledRed          : out   slv(1 downto 0);
      ledGrn          : out   slv(1 downto 0);
      ledBlu          : out   slv(1 downto 0);
      -- Stable Reference IDELAY Clock and Reset
      refClk200MHz    : in    sl;
      refRst200MHz    : in    sl;
      -- Camera Control Bits
      camCtrl         : in    Slv4Array(1 downto 0);
      -- Camera Data Interface
      dataMasters     : out   AxiStreamMasterArray(1 downto 0) := (others => AXI_STREAM_MASTER_INIT_C);
      dataSlaves      : in    AxiStreamSlaveArray(1 downto 0);
      -- UART Interface
      rxUartMasters   : in    AxiStreamMasterArray(1 downto 0);
      rxUartSlaves    : out   AxiStreamSlaveArray(1 downto 0)  := (others => AXI_STREAM_SLAVE_FORCE_C);
      txUartMasters   : out   AxiStreamMasterArray(1 downto 0) := (others => AXI_STREAM_MASTER_INIT_C);
      txUartSlaves    : in    AxiStreamSlaveArray(1 downto 0);
      -- Axi-Lite Interface
      axilClk         : in    sl;
      axilRst         : in    sl;
      axilReadMaster  : in    AxiLiteReadMasterType;
      axilReadSlave   : out   AxiLiteReadSlaveType;
      axilWriteMaster : in    AxiLiteWriteMasterType;
      axilWriteSlave  : out   AxiLiteWriteSlaveType);
end CLinkWrapper;

architecture mapping of CLinkWrapper is

   signal txMasterA : AxiStreamMasterArray(CHAN_COUNT_G-1 downto 0);
   signal txSlaveA  : AxiStreamSlaveArray(CHAN_COUNT_G-1 downto 0);

   signal txMasterB : AxiStreamMasterArray(CHAN_COUNT_G-1 downto 0);
   signal txSlaveB  : AxiStreamSlaveArray(CHAN_COUNT_G-1 downto 0);

   signal txMasterC : AxiStreamMasterArray(CHAN_COUNT_G-1 downto 0);
   signal txSlaveC  : AxiStreamSlaveArray(CHAN_COUNT_G-1 downto 0);

   signal camStatus : ClChanStatusArray(1 downto 0);

begin

   U_ClinkTop : entity surf.ClinkTop
      generic map (
         TPD_G              => TPD_G,
         CHAN_COUNT_G       => CHAN_COUNT_G,
         UART_READY_EN_G    => true,
         COMMON_AXIL_CLK_G  => true,
         COMMON_DATA_CLK_G  => true,
         DATA_AXIS_CONFIG_G => PGP3_AXIS_CONFIG_C,
         UART_AXIS_CONFIG_G => PGP3_AXIS_CONFIG_C,
         AXIL_BASE_ADDR_G   => AXIL_BASE_ADDR_G)
      port map (
         -- Clink Ports
         cbl0Half0P      => cbl0Half0P,
         cbl0Half0M      => cbl0Half0M,
         cbl0Half1P      => cbl0Half1P,
         cbl0Half1M      => cbl0Half1M,
         cbl0SerP        => cbl0SerP,
         cbl0SerM        => cbl0SerM,
         cbl1Half0P      => cbl1Half0P,
         cbl1Half0M      => cbl1Half0M,
         cbl1Half1P      => cbl1Half1P,
         cbl1Half1M      => cbl1Half1M,
         cbl1SerP        => cbl1SerP,
         cbl1SerM        => cbl1SerM,
         -- Delay clock and reset, 200Mhz
         dlyClk          => refClk200MHz,
         dlyRst          => refRst200MHz,
         -- System clock and reset, > 100 Mhz
         sysClk          => axilClk,
         sysRst          => axilRst,
         -- Camera Control Bits & status, async
         camCtrl         => camCtrl(CHAN_COUNT_G-1 downto 0),
         camStatus       => camStatus,
         -- Camera data
         dataClk         => axilClk,
         dataRst         => axilRst,
         dataMasters     => dataMasters(CHAN_COUNT_G-1 downto 0),
         dataSlaves      => dataSlaves(CHAN_COUNT_G-1 downto 0),
         -- UART data
         uartClk         => axilClk,
         uartRst         => axilRst,
         sUartMasters    => rxUartMasters(CHAN_COUNT_G-1 downto 0),
         sUartSlaves     => rxUartSlaves(CHAN_COUNT_G-1 downto 0),
         mUartMasters    => txUartMasters(CHAN_COUNT_G-1 downto 0),
         mUartSlaves     => txUartSlaves(CHAN_COUNT_G-1 downto 0),
         -- Axi-Lite Interface
         axilClk         => axilClk,
         axilRst         => axilRst,
         axilReadMaster  => axilReadMaster,
         axilReadSlave   => axilReadSlave,
         axilWriteMaster => axilWriteMaster,
         axilWriteSlave  => axilWriteSlave);

   ----------------
   -- Misc. Signals
   ----------------
   process (camStatus)
   begin

      if camStatus(0).running = '1' then
         ledRed(0) <= '1';
         ledGrn(0) <= '0';
         ledBlu(0) <= '1';
      else
         ledRed(0) <= '0';
         ledGrn(0) <= '1';
         ledBlu(0) <= '1';
      end if;

      if CHAN_COUNT_G = 1 then
         ledRed(1) <= '1';
         ledGrn(1) <= '1';
         ledBlu(1) <= '1';
      elsif camStatus(1).running = '1' then
         ledRed(1) <= '1';
         ledGrn(1) <= '0';
         ledBlu(1) <= '1';
      else
         ledRed(1) <= '0';
         ledGrn(1) <= '1';
         ledBlu(1) <= '1';
      end if;

   end process;

end mapping;
